`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    20:08:50 10/09/2019 
// Design Name: 
// Module Name:    location_judge 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module location_judge(
    clk,rst_n,save_en,fetch_en,location_coding,rotate_direction,rotate_en,rise_fall_direction,rise_fall_en,rise_fall_en_main,
	extend_shrink_direction,extend_shrink_en,occupy_en,empty_location_en,accomplish_en,yuyin_end_en
	);
	input clk;
	input rst_n;
	input save_en;    //存储信号
	input fetch_en;      //取物信号
	input [6:0] location_coding;   //位置编码(seven)
	
	output  reg occupy_en;      //工作信号（高电平表示正在工作）   occupy（vi占据，占领，居住，使忙碌）
	output  reg empty_location_en;    //清空地址，使能信号（高电平时对地址进行清零）
	output  reg accomplish_en;    //完成信号
	
	output  reg rotate_direction;   //旋转方向信号（0：顺时针；1：逆时针）
	output  reg rotate_en;   //旋转使能信号
	output  reg rise_fall_direction;   //升降方向信号（0：上升；1：下降）
	output  reg rise_fall_en;     //升降使能信号
	output  reg rise_fall_en_main;    //大幅度升降使能信号
	output  reg extend_shrink_direction;  //伸缩方向信号（0：伸长；1：缩回）
	output	reg extend_shrink_en;   //伸缩使能信号
	output reg [1:0]yuyin_end_en;
	reg [31:0]rotate_cnt;   //旋转数值
	reg [31:0]rise_fall_cnt;   //升降数值
	reg [31:0]extend_shrink_cnt;     //伸缩数值
	
	reg [31:0]cnt_c;   //旋转计数器
	reg [31:0]cnt_b;   //升降计数器
	reg [31:0]cnt_a;     //伸缩计数器
	
	reg extend_shrink_end;   //伸缩停止信号(高电平有效)
	reg rise_fall_end;        //升降停止信号(高电平有效)
	reg rotate_end;           //旋转停止信号(高电平有效)
	
	reg reset_cnt;   //计数器清零信号
	
/* 	parameter  ROTATE_CNT_A=32'd8000 ,     //旋转角度固定值
	           ROTATE_CNT_B=32'd8000 ;    
	parameter RISE_FALL_CNT_A=32'd6000,    //升降距离固定值
	          RISE_FALL_CNT_B=32'd1000 ;
	parameter  EXTEND_SHRINK_CNT_A=32'd7000,    //伸缩长度固定值
	           EXTEND_SHRINK_CNT_B=32'd7000;
	 */		   
	parameter  ROTATE_CNT_A=32'd24_000_000*4'd3+32'd15_000_000 ,     //旋转角度固定值
	           ROTATE_CNT_B=32'd24_000_000 ;    
	parameter RISE_FALL_CNT_A=32'd24_000_000*4'd6+32'd19_000_000,    //升降距离固定值
	          RISE_FALL_CNT_B=32'd24_000_000*4'd4 ;
	parameter  EXTEND_SHRINK_CNT_A=32'd24_000_000*4'd5+32'd16_000_000,    //伸缩长度固定值
	           EXTEND_SHRINK_CNT_B=32'd24_000_000*4'd5+32'd16_000_000; 
	
	reg [6:0]current_state;   //现态
	reg [6:0]next_state;    //下一个状态
	reg [6:0]last_state;   //上一个状态
	
	parameter   S0=7'b000_000_0,S1=7'b000_000_1,S2=7'b001_000_1,S3=7'b001_000_0,        //初始位置
	            
				AQ1=7'b000_001_0,AQ2=7'b000_001_1,AQ3=7'b001_001_1,AQ4=7'b001_001_0,    //第一层
				AW1=7'b000_010_0,AW2=7'b000_010_1,AW3=7'b001_010_1,AW4=7'b001_010_0,
				AE1=7'b000_011_0,AE2=7'b000_011_1,AE3=7'b001_011_1,AE4=7'b001_011_0,
				AR1=7'b000_100_0,AR2=7'b000_100_1,AR3=7'b001_100_1,AR4=7'b001_100_0,
				
				BQ1=7'b010_001_0,BQ2=7'b010_001_1,BQ3=7'b011_001_1,BQ4=7'b011_001_0,    //第二层
				BW1=7'b010_010_0,BW2=7'b010_010_1,BW3=7'b011_010_1,BW4=7'b011_010_0,
				BE1=7'b010_011_0,BE2=7'b010_011_1,BE3=7'b011_011_1,BE4=7'b011_011_0,
				BR1=7'b010_100_0,BR2=7'b010_100_1,BR3=7'b011_100_1,BR4=7'b011_100_0,
				
				CQ1=7'b100_001_0,CQ2=7'b100_001_1,CQ3=7'b101_001_1,CQ4=7'b101_001_0,    //第三层
				CW1=7'b100_010_0,CW2=7'b100_010_1,CW3=7'b101_010_1,CW4=7'b101_010_0,
				CE1=7'b100_011_0,CE2=7'b100_011_1,CE3=7'b101_011_1,CE4=7'b101_011_0,
				CR1=7'b100_100_0,CR2=7'b100_100_1,CR3=7'b101_100_1,CR4=7'b101_100_0,
				
				DQ1=7'b110_001_0,DQ2=7'b110_001_1,DQ3=7'b111_001_1,DQ4=7'b111_001_0,     //第四层
				DW1=7'b110_010_0,DW2=7'b110_010_1,DW3=7'b111_010_1,DW4=7'b111_010_0,
				DE1=7'b110_011_0,DE2=7'b110_011_1,DE3=7'b111_011_1,DE4=7'b111_011_0,
				DR1=7'b110_100_0,DR2=7'b110_100_1,DR3=7'b111_100_1,DR4=7'b111_100_0;
	
	always@(posedge clk or negedge rst_n)
	begin
	if(!rst_n)
		begin
		current_state<=7'd0;
		end
	else
		begin
		current_state<=next_state;
		end
	end
	
	always@(posedge clk or negedge rst_n)
	begin
	if(!rst_n)
	begin
	occupy_en<=1'b0;
	rotate_en<=1'b0;
	rotate_direction<=1'b0;
	rotate_cnt<=32'd0;
	extend_shrink_en<=1'b0;
	extend_shrink_cnt<=32'd0;
	extend_shrink_direction<=1'b0;
	rise_fall_en<=1'b0;
	rise_fall_en_main<=1'b0;
	rise_fall_cnt<=32'd0;     
	rise_fall_direction<=1'b0;
	accomplish_en<=1'b0;
	reset_cnt<=1'b1;
	yuyin_end_en<=2'b00;
	end
	else
		begin
		case(current_state)
		S0:begin
			empty_location_en<=1'b0;
		    if(save_en)             
		    begin
				accomplish_en<=1'b0;
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b0;
				yuyin_end_en<=2'b00;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;     
			    if(!extend_shrink_end)
			        begin
					next_state<=S0;
			    	end
			    else
					begin
					next_state<=S1;
					last_state<=S0;
			    	end
			end
			else if(fetch_en)
			    begin
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b1;
				extend_shrink_cnt<=(EXTEND_SHRINK_CNT_A*(last_state[0]-current_state[0]));
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=S0;
					occupy_en<=1'b1;
					yuyin_end_en<=2'b00;
					accomplish_en<=1'b0;
			    	end
			    else
					begin
					next_state<=location_coding;
					occupy_en<=1'b0;
					accomplish_en<=1'b1;
					yuyin_end_en<=2'b00;
					last_state<=S0;
			    	end
				end
			else
				begin
				yuyin_end_en<=2'b00;
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				accomplish_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=S0;
				end
		   end
		S1:begin
			accomplish_en<=1'b0;
			empty_location_en<=1'b0;
			if(save_en)
				begin
				yuyin_end_en<=2'b00;
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b0;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b1;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=RISE_FALL_CNT_B;     
			    rise_fall_direction<=1'b0;	
				if(!rise_fall_end)
			        begin
					next_state<=S1;
			    	end
			    else
					begin
					next_state<=S2;
					last_state<=S1;
			    	end
				end
			else if(fetch_en)
				begin
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b0;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b1;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=RISE_FALL_CNT_B;     
			    rise_fall_direction<=1'b1;	
				if(!rise_fall_end)
			        begin
					next_state<=S1;
					yuyin_end_en<=2'b00;
			    	end
			    else
					begin
					next_state<=S0;
					last_state<=S1;
					yuyin_end_en<=2'b10;
			    	end
				end
			else
				begin
				yuyin_end_en<=2'b00;
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=S1;
				end
		   end
		S2:begin
			empty_location_en<=1'b0;
			yuyin_end_en<=2'b00;
			accomplish_en<=1'b0;
			if(save_en)
				begin
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b1;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=S2;
			    	end
			    else
					begin
					last_state<=S2;
					next_state<=S3;
			    	end
				end
			else if(fetch_en)
				begin
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;     //伸缩长度
			    if(!extend_shrink_end)
			        begin
					next_state<=S2;
			    	end
			    else
					begin
					last_state<=S2;
					next_state<=S1;
			    	end
			    end
			else
				begin
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=S2;
				end
		   end
		S3:begin
			yuyin_end_en<=2'b00;
			accomplish_en<=1'b0;
			if(save_en)
				begin
				occupy_en<=1'b1;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b0;
				if(!rise_fall_end)
					begin
					rise_fall_en_main<=1'b1;
					end
				else
					begin
					rise_fall_en_main<=1'b0;
					end
				if(!rotate_end)
					begin
					rotate_en<=1'b1;
					end
				else
					begin
					rotate_en<=1'b0;
					end
					
				if(location_coding[6:5]>current_state[6:5])
					begin
					rise_fall_cnt<=(location_coding[6:5]-current_state[6:5])*RISE_FALL_CNT_A;     //升的高度
					rise_fall_direction<=1'b0;
					end
				else
					begin
					rise_fall_cnt<=(current_state[6:5]-location_coding[6:5])*RISE_FALL_CNT_A;     //降的高度
					rise_fall_direction<=1'b1;
					end
				if(location_coding[3:1]>current_state[3:1])
				    begin
				    rotate_cnt<=(location_coding[3:1]-current_state[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b0;
				    end
				else
				    begin
				    rotate_cnt<=(current_state[3:1]-location_coding[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b1;
				    end
				
			    if((!rise_fall_end)|(!rotate_end))
				    begin
					next_state<=S3;
					empty_location_en<=1'b0;
					reset_cnt<=1'b0;
				    end
				else
					begin
					last_state<=S3;
					empty_location_en<=1'b1;
					next_state<=location_coding;
					reset_cnt<=1'b1;
					end
			
		        end
			else if(fetch_en)
				begin
				occupy_en<=1'b1;
				empty_location_en<=1'b0;
				
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b0;
				if(!rise_fall_end)
					begin
					rise_fall_en_main<=1'b1;
					end
				else
					begin
					rise_fall_en_main<=1'b0;
					end
				if(!rotate_end)
					begin
					rotate_en<=1'b1;
					end
				else
					begin
					rotate_en<=1'b0;
					end
					
				
				if(last_state[6:5]>current_state[6:5])
					begin
					rise_fall_cnt<=(last_state[6:5]-current_state[6:5])*RISE_FALL_CNT_A;     //升的高度
					rise_fall_direction<=1'b1;
					end
				else
					begin
					rise_fall_cnt<=(current_state[6:5]-last_state[6:5])*RISE_FALL_CNT_A;     //降的高度
					rise_fall_direction<=1'b0;
					end
				if(last_state[3:1]>current_state[3:1])
				    begin
				    rotate_cnt<=(last_state[3:1]-current_state[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b1;
				    end
				else
				    begin
				    rotate_cnt<=(current_state[3:1]-last_state[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b0;
				    end
			    if((!rise_fall_end)|(!rotate_end))
				    begin
					next_state<=S3;
					reset_cnt<=1'b0;
				    end
				else
					begin
					next_state<=S2;
					last_state<=S3;
					reset_cnt<=1'b1;
					end
			    end
		        
			else
				begin
				occupy_en<=1'b0;
				empty_location_en<=1'b0;
				
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=S3;
				end
		   end
		   
//第一层	
		//第一层顺时针第一个房间
		AQ1:begin
			accomplish_en<=1'b0;
			yuyin_end_en<=2'b00;
		    if(fetch_en)
		    begin
				occupy_en<=1'b1;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b0;
				if(!rise_fall_end)
					begin
					rise_fall_en_main<=1'b1;
					end
				else
					begin
					rise_fall_en_main<=1'b0;
					end
				if(!rotate_end)
					begin
					rotate_en<=1'b1;
					end
				else
					begin
					rotate_en<=1'b0;
					end
					
				if(location_coding[6:5]>last_state[6:5])
					begin
					rise_fall_cnt<=(location_coding[6:5]-last_state[6:5])*RISE_FALL_CNT_A;     //升的高度
					rise_fall_direction<=1'b0;
					end
				else
					begin
					rise_fall_cnt<=(last_state[6:5]-location_coding[6:5])*RISE_FALL_CNT_A;     //降的高度
					rise_fall_direction<=1'b1;
					end
				if(location_coding[3:1]>last_state[3:1])
				    begin
				    rotate_cnt<=(location_coding[3:1]-last_state[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b0;
				    end
				else
				    begin
				    rotate_cnt<=(last_state[3:1]-location_coding[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b1;
				    end
			    if((!rise_fall_end)|(!rotate_end))
				    begin
					next_state<=AQ1;
					reset_cnt<=1'b0;
				    end
				else
					begin
					next_state<={location_coding[6:1],1'b1};
					empty_location_en<=1'b1;
					last_state<=AQ1;
					reset_cnt<=1'b1;
					end
			
		    end
			else if(save_en)
			    begin
				occupy_en<=1'b1;
				empty_location_en<=1'b0;
				
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b0;
				if(!rise_fall_end)
					begin
					rise_fall_en_main<=1'b1;
					end
				else
					begin
					rise_fall_en_main<=1'b0;
					end
				if(!rotate_end)
					begin
					rotate_en<=1'b1;
					end
				else
					begin
					rotate_en<=1'b0;
					end
					
				if(S0[6:5]>current_state[6:5])
					begin
					rise_fall_cnt<=(S0[6:5]-current_state[6:5])*RISE_FALL_CNT_A;     //升的高度
					rise_fall_direction<=1'b0;
					end
				else
					begin
					rise_fall_cnt<=(current_state[6:5]-S0[6:5])*RISE_FALL_CNT_A;     //降的高度
					rise_fall_direction<=1'b1;
					end
				if(S0[3:1]>current_state[3:1])
				    begin
				    rotate_cnt<=(S0[3:1]-current_state[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b0;
				    end
				else
				    begin
				    rotate_cnt<=(current_state[3:1]-S0[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b1;
				    end
			    if((!rise_fall_end)|(!rotate_end))
				    begin
					next_state<=AQ1;
					reset_cnt<=1'b0;
					
				    end
				else
					begin
					next_state<=S0;
					last_state<=AQ1;
					reset_cnt<=1'b1;
					end
			
		        end
			else
				begin
				empty_location_en<=1'b0;
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=AQ1;
				end
		   end
		AQ2:begin
			empty_location_en<=1'b0;
			if(fetch_en)
				begin
				yuyin_end_en<=2'b00;
				accomplish_en<=1'b0;
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=AQ2;
			    	end
			    else
					begin
					last_state<=AQ2;
					next_state<=AQ3;
			    	end
				end
			else if(save_en)
				begin
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b1;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=AQ2;
					occupy_en<=1'b1;
					yuyin_end_en<=2'b00;
					accomplish_en<=1'b0;
			    	end
			    else
					begin
					last_state<=AQ2;
					next_state<=AQ1;
					occupy_en<=1'b0;
					yuyin_end_en<=2'b01;
					accomplish_en<=1'b1;
			    	end
				end
			else
				begin
				occupy_en<=1'b0;
				accomplish_en<=1'b0;
				rotate_en<=1'b0;
				yuyin_end_en<=2'b00;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=AQ2;
				end
		   end
		AQ3:begin
			empty_location_en<=1'b0;
			yuyin_end_en<=2'b00;
			if(fetch_en)
				begin
				occupy_en<=1'b1;
				
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b0;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b1;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=RISE_FALL_CNT_B;     
			    rise_fall_direction<=1'b0;	
				if(!rise_fall_end)
			        begin
					next_state<=AQ3;
			    	end
			    else
					begin
					last_state<=AQ3;
					next_state<=AQ4;
			    	end
				end
			else if(save_en)
				begin
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b0;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b1;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=RISE_FALL_CNT_B;     
			    rise_fall_direction<=1'b1;	
				if(!rise_fall_end)
			        begin
					next_state<=AQ3;
			    	end
			    else
					begin
					last_state<=AQ3;
					next_state<=AQ2;
			    	end
				end
			else
				begin
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=AQ3;
				end
		   end
		AQ4:begin
			empty_location_en<=1'b0;
			yuyin_end_en<=2'b00;
			if(fetch_en)
				begin
				occupy_en<=1'b1;
				
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b1;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=AQ4;
			    	end
			    else
					begin
					last_state<=AQ4;
					next_state<=S3;
			    	end
				end
			else if(save_en)
				begin
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;     //伸缩长度
			    if(!extend_shrink_end)
			        begin
					next_state<=AQ4;
			    	end
			    else
					begin
					last_state<=AQ4;
					next_state<=AQ3;
			    	end
			    end
			else
				begin
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=AQ4;
				end
		   end
		//第一层顺时针第二个房间 
		AW1:begin
			accomplish_en<=1'b0;
			yuyin_end_en<=2'b00;
		    if(fetch_en)
		    begin
				occupy_en<=1'b1;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b0;
				if(!rise_fall_end)
					begin
					rise_fall_en_main<=1'b1;
					end
				else
					begin
					rise_fall_en_main<=1'b0;
					end
				if(!rotate_end)
					begin
					rotate_en<=1'b1;
					end
				else
					begin
					rotate_en<=1'b0;
					end
					
				if(location_coding[6:5]>last_state[6:5])
					begin
					rise_fall_cnt<=(location_coding[6:5]-last_state[6:5])*RISE_FALL_CNT_A;     //升的高度
					rise_fall_direction<=1'b0;
					end
				else
					begin
					rise_fall_cnt<=(last_state[6:5]-location_coding[6:5])*RISE_FALL_CNT_A;     //降的高度
					rise_fall_direction<=1'b1;
					end
				if(location_coding[3:1]>last_state[3:1])
				    begin
				    rotate_cnt<=(location_coding[3:1]-last_state[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b0;
				    end
				else
				    begin
				    rotate_cnt<=(last_state[3:1]-location_coding[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b1;
				    end
			    if((!rise_fall_end)|(!rotate_end))
				    begin
					next_state<=AW1;
					reset_cnt<=1'b0;
				    end
				else
					begin
					reset_cnt<=1'b1;
					next_state<={location_coding[6:1],1'b1};
					empty_location_en<=1'b1;
					last_state<=AW1;
					end
			
		    end
			else if(save_en)
			    begin
				occupy_en<=1'b1;
				empty_location_en<=1'b0;
				
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b0;
				if(!rise_fall_end)
					begin
					rise_fall_en_main<=1'b1;
					end
				else
					begin
					rise_fall_en_main<=1'b0;
					end
				if(!rotate_end)
					begin
					rotate_en<=1'b1;
					end
				else
					begin
					rotate_en<=1'b0;
					end
					
				if(S0[6:5]>current_state[6:5])
					begin
					rise_fall_cnt<=(S0[6:5]-current_state[6:5])*RISE_FALL_CNT_A;     //升的高度
					rise_fall_direction<=1'b0;
					end
				else
					begin
					rise_fall_cnt<=(current_state[6:5]-S0[6:5])*RISE_FALL_CNT_A;     //降的高度
					rise_fall_direction<=1'b1;
					end
				if(S0[3:1]>current_state[3:1])
				    begin
				    rotate_cnt<=(S0[3:1]-current_state[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b0;
				    end
				else
				    begin
				    rotate_cnt<=(current_state[3:1]-S0[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b1;
				    end
			    if((!rise_fall_end)|(!rotate_end))
				    begin
					next_state<=AW1;
					reset_cnt<=1'b0;
				    end
				else
					begin
					next_state<=S0;
					last_state<=AW1;
					reset_cnt<=1'b1;
					end
			
		        end
			else
				begin
				empty_location_en<=1'b0;
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=AW1;
				end
		   end
		AW2:begin
			empty_location_en<=1'b0;
			if(fetch_en)
				begin
				yuyin_end_en<=2'b00;
				accomplish_en<=1'b0;
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=AW2;
			    	end
			    else
					begin
					last_state<=AW2;
					next_state<=AW3;
			    	end
				end
			else if(save_en)
				begin
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b1;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=AW2;
					occupy_en<=1'b1;
					accomplish_en<=1'b0;
					yuyin_end_en<=2'b00;
			    	end
			    else
					begin
					last_state<=AW2;
					next_state<=AW1;
					occupy_en<=1'b0;
					accomplish_en<=1'b1;
					yuyin_end_en<=2'b01;
			    	end
				end
			else
				begin
				yuyin_end_en<=2'b00;
				occupy_en<=1'b0;
				accomplish_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=AW2;
				end
		   end
		AW3:begin
			empty_location_en<=1'b0;
			yuyin_end_en<=2'b00;
			if(fetch_en)
				begin
				occupy_en<=1'b1;
				
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b0;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b1;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=RISE_FALL_CNT_B;     
			    rise_fall_direction<=1'b0;	
				if(!rise_fall_end)
			        begin
					next_state<=AW3;
			    	end
			    else
					begin
					last_state<=AW3;
					next_state<=AW4;
			    	end
				end
			else if(save_en)
				begin
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b0;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b1;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=RISE_FALL_CNT_B;     
			    rise_fall_direction<=1'b1;	
				if(!rise_fall_end)
			        begin
					next_state<=AW3;
			    	end
			    else
					begin
					last_state<=AW3;
					next_state<=AW2;
			    	end
				end
			else
				begin
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=AW3;
				end
		   end
		AW4:begin
			empty_location_en<=1'b0;
			yuyin_end_en<=2'b00;
			if(fetch_en)
				begin
				occupy_en<=1'b1;
				
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b1;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=AW4;
			    	end
			    else
					begin
					last_state<=AW4;
					next_state<=S3;
			    	end
				end
			else if(save_en)
				begin
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;     //伸缩长度
			    if(!extend_shrink_end)
			        begin
					next_state<=AW4;
			    	end
			    else
					begin
					last_state<=AW4;
					next_state<=AW3;
			    	end
			    end
			else
				begin
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=AW4;
				end
		   end
		//第一层顺时针第三个房间
		AE1:begin
			accomplish_en<=1'b0;
			yuyin_end_en<=2'b00;
		    if(fetch_en)
		    begin
				occupy_en<=1'b1;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b0;
				if(!rise_fall_end)
					begin
					rise_fall_en_main<=1'b1;
					end
				else
					begin
					rise_fall_en_main<=1'b0;
					end
				if(!rotate_end)
					begin
					rotate_en<=1'b1;
					end
				else
					begin
					rotate_en<=1'b0;
					end
					
				if(location_coding[6:5]>last_state[6:5])
					begin
					rise_fall_cnt<=(location_coding[6:5]-last_state[6:5])*RISE_FALL_CNT_A;     //升的高度
					rise_fall_direction<=1'b0;
					end
				else
					begin
					rise_fall_cnt<=(last_state[6:5]-location_coding[6:5])*RISE_FALL_CNT_A;     //降的高度
					rise_fall_direction<=1'b1;
					end
				if(location_coding[3:1]>last_state[3:1])
				    begin
				    rotate_cnt<=(location_coding[3:1]-last_state[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b0;
				    end
				else
				    begin
				    rotate_cnt<=(last_state[3:1]-location_coding[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b1;
				    end
			    if((!rise_fall_end)|(!rotate_end))
				    begin
					next_state<=AE1;
					reset_cnt<=1'b0;
				    end
				else
					begin
					reset_cnt<=1'b1;
					next_state<={location_coding[6:1],1'b1};
					empty_location_en<=1'b1;
					last_state<=AE1;
					end
			
		    end
			else if(save_en)
			    begin
				occupy_en<=1'b1;
				empty_location_en<=1'b0;
				
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b0;
				if(!rise_fall_end)
					begin
					rise_fall_en_main<=1'b1;
					end
				else
					begin
					rise_fall_en_main<=1'b0;
					end
				if(!rotate_end)
					begin
					rotate_en<=1'b1;
					end
				else
					begin
					rotate_en<=1'b0;
					end
					
				if(S0[6:5]>current_state[6:5])
					begin
					rise_fall_cnt<=(S0[6:5]-current_state[6:5])*RISE_FALL_CNT_A;     //升的高度
					rise_fall_direction<=1'b0;
					end
				else
					begin
					rise_fall_cnt<=(current_state[6:5]-S0[6:5])*RISE_FALL_CNT_A;     //降的高度
					rise_fall_direction<=1'b1;
					end
				if(S0[3:1]>current_state[3:1])
				    begin
				    rotate_cnt<=(S0[3:1]-current_state[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b0;
				    end
				else
				    begin
				    rotate_cnt<=(current_state[3:1]-S0[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b1;
				    end
			    if((!rise_fall_end)|(!rotate_end))
				    begin
					next_state<=AE1;
					reset_cnt<=1'b0;
				    end
				else
					begin
					next_state<=S0;
					last_state<=AE1;
					reset_cnt<=1'b1;
					end
			
		        end
			else
				begin
				empty_location_en<=1'b0;
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=AE1;
				end
		   end
		AE2:begin
			empty_location_en<=1'b0;
			if(fetch_en)
				begin
				yuyin_end_en<=2'b00;
				accomplish_en<=1'b0;
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=AE2;
			    	end
			    else
					begin
					last_state<=AE2;
					next_state<=AE3;
			    	end
				end
			else if(save_en)
				begin
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b1;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=AE2;
					occupy_en<=1'b1;
					yuyin_end_en<=2'b00;
					accomplish_en<=1'b0;
			    	end
			    else
					begin
					last_state<=AE2;
					next_state<=AE1;
					occupy_en<=1'b0;
					yuyin_end_en<=2'b01;
					accomplish_en<=1'b1;
			    	end
				end
			else
				begin
				yuyin_end_en<=2'b00;
				occupy_en<=1'b0;
				accomplish_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=AE2;
				end
		   end
		AE3:begin
			empty_location_en<=1'b0;
			yuyin_end_en<=2'b00;
			if(fetch_en)
				begin
				occupy_en<=1'b1;
				
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b0;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b1;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=RISE_FALL_CNT_B;     
			    rise_fall_direction<=1'b0;	
				if(!rise_fall_end)
			        begin
					next_state<=AE3;
			    	end
			    else
					begin
					last_state<=AE3;
					next_state<=AE4;
			    	end
				end
			else if(save_en)
				begin
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b0;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b1;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=RISE_FALL_CNT_B;     
			    rise_fall_direction<=1'b1;	
				if(!rise_fall_end)
			        begin
					next_state<=AE3;
			    	end
			    else
					begin
					last_state<=AE3;
					next_state<=AE2;
			    	end
				end
			else
				begin
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=AE3;
				end
		   end
		AE4:begin
			empty_location_en<=1'b0;
			yuyin_end_en<=2'b00;
			if(fetch_en)
				begin
				occupy_en<=1'b1;
				
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b1;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=AE4;
			    	end
			    else
					begin
					last_state<=AE4;
					next_state<=S3;
			    	end
				end
			else if(save_en)
				begin
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;     //伸缩长度
			    if(!extend_shrink_end)
			        begin
					next_state<=AE4;
			    	end
			    else
					begin
					last_state<=AE4;
					next_state<=AE3;
			    	end
			    end
			else
				begin
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=AE4;
				end
		   end
		//第一层顺时针第四个房间
		AR1:begin
			accomplish_en<=1'b0;
			yuyin_end_en<=2'b00;
		    if(fetch_en)
		    begin
				occupy_en<=1'b1;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b0;
				if(!rise_fall_end)
					begin
					rise_fall_en_main<=1'b1;
					end
				else
					begin
					rise_fall_en_main<=1'b0;
					end
				if(!rotate_end)
					begin
					rotate_en<=1'b1;
					end
				else
					begin
					rotate_en<=1'b0;
					end
					
				if(location_coding[6:5]>last_state[6:5])
					begin
					rise_fall_cnt<=(location_coding[6:5]-last_state[6:5])*RISE_FALL_CNT_A;     //升的高度
					rise_fall_direction<=1'b0;
					end
				else
					begin
					rise_fall_cnt<=(last_state[6:5]-location_coding[6:5])*RISE_FALL_CNT_A;     //降的高度
					rise_fall_direction<=1'b1;
					end
				if(location_coding[3:1]>last_state[3:1])
				    begin
				    rotate_cnt<=(location_coding[3:1]-last_state[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b0;
				    end
				else
				    begin
				    rotate_cnt<=(last_state[3:1]-location_coding[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b1;
				    end
			    if((!rise_fall_end)|(!rotate_end))
				    begin
					next_state<=AR1;
					reset_cnt<=1'b0;
				    end
				else
					begin
					next_state<={location_coding[6:1],1'b1};
					empty_location_en<=1'b1;
					last_state<=AR1;
					reset_cnt<=1'b1;
					end
			
		    end
			else if(save_en)
			    begin
				occupy_en<=1'b1;
				empty_location_en<=1'b0;
				
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b0;
				if(!rise_fall_end)
					begin
					rise_fall_en_main<=1'b1;
					end
				else
					begin
					rise_fall_en_main<=1'b0;
					end
				if(!rotate_end)
					begin
					rotate_en<=1'b1;
					end
				else
					begin
					rotate_en<=1'b0;
					end
					
				if(S0[6:5]>current_state[6:5])
					begin
					rise_fall_cnt<=(S0[6:5]-current_state[6:5])*RISE_FALL_CNT_A;     //升的高度
					rise_fall_direction<=1'b0;
					end
				else
					begin
					rise_fall_cnt<=(current_state[6:5]-S0[6:5])*RISE_FALL_CNT_A;     //降的高度
					rise_fall_direction<=1'b1;
					end
				if(S0[3:1]>current_state[3:1])
				    begin
				    rotate_cnt<=(S0[3:1]-current_state[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b0;
				    end
				else
				    begin
				    rotate_cnt<=(current_state[3:1]-S0[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b1;
				    end
			    if((!rise_fall_end)|(!rotate_end))
				    begin
					next_state<=AR1;
					reset_cnt<=1'b0;
				    end
				else
					begin
					next_state<=S0;
					last_state<=AR1;
					reset_cnt<=1'b1;
					end
			
		        end
			else
				begin
				empty_location_en<=1'b0;
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=AR1;
				end
		   end
		AR2:begin
			empty_location_en<=1'b0;
			if(fetch_en)
				begin
				yuyin_end_en<=2'b00;
				accomplish_en<=1'b0;
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=AR2;
			    	end
			    else
					begin
					last_state<=AR2;
					next_state<=AR3;
			    	end
				end
			else if(save_en)
				begin
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b1;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=AR2;
					occupy_en<=1'b1;
					yuyin_end_en<=2'b00;
					accomplish_en<=1'b0;
			    	end
			    else
					begin
					last_state<=AR2;
					next_state<=AR1;
					occupy_en<=1'b0;
					yuyin_end_en<=2'b01;
					accomplish_en<=1'b1;
			    	end
				end
			else
				begin
				yuyin_end_en<=2'b00;
				accomplish_en<=1'b0;
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=AR2;
				end
		   end
		AR3:begin
			empty_location_en<=1'b0;
			yuyin_end_en<=2'b00;
			if(fetch_en)
				begin
				occupy_en<=1'b1;
				
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b0;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b1;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=RISE_FALL_CNT_B;     
			    rise_fall_direction<=1'b0;	
				if(!rise_fall_end)
			        begin
					next_state<=AR3;
			    	end
			    else
					begin
					last_state<=AR3;
					next_state<=AR4;
			    	end
				end
			else if(save_en)
				begin
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b0;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b1;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=RISE_FALL_CNT_B;     
			    rise_fall_direction<=1'b1;	
				if(!rise_fall_end)
			        begin
					next_state<=AR3;
			    	end
			    else
					begin
					last_state<=AR3;
					next_state<=AR2;
			    	end
				end
			else
				begin
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=AR3;
				end
		   end
		AR4:begin
			empty_location_en<=1'b0;
			yuyin_end_en<=2'b00;
			if(fetch_en)
				begin
				occupy_en<=1'b1;
				
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b1;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=AR4;
			    	end
			    else
					begin
					last_state<=AR4;
					next_state<=S3;
			    	end
				end
			else if(save_en)
				begin
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;     //伸缩长度
			    if(!extend_shrink_end)
			        begin
					next_state<=AR4;
			    	end
			    else
					begin
					last_state<=AR4;
					next_state<=AR3;
			    	end
			    end
			else
				begin
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=AR4;
				end
		   end
		
//第二层
		//第二层顺时针第一个房间
        BQ1:begin
			accomplish_en<=1'b0;
			yuyin_end_en<=2'b00;
		    if(fetch_en)
		    begin
				occupy_en<=1'b1;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b0;
				if(!rise_fall_end)
					begin
					rise_fall_en_main<=1'b1;
					end
				else
					begin
					rise_fall_en_main<=1'b0;
					end
				if(!rotate_end)
					begin
					rotate_en<=1'b1;
					end
				else
					begin
					rotate_en<=1'b0;
					end
					
				if(location_coding[6:5]>last_state[6:5])
					begin
					rise_fall_cnt<=(location_coding[6:5]-last_state[6:5])*RISE_FALL_CNT_A;     //升的高度
					rise_fall_direction<=1'b0;
					end
				else
					begin
					rise_fall_cnt<=(last_state[6:5]-location_coding[6:5])*RISE_FALL_CNT_A;     //降的高度
					rise_fall_direction<=1'b1;
					end
				if(location_coding[3:1]>last_state[3:1])
				    begin
				    rotate_cnt<=(location_coding[3:1]-last_state[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b0;
				    end
				else
				    begin
				    rotate_cnt<=(last_state[3:1]-location_coding[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b1;
				    end
			    if((!rise_fall_end)|(!rotate_end))
				    begin
					next_state<=BQ1;
					reset_cnt<=1'b0;
				    end
				else
					begin
					next_state<={location_coding[6:1],1'b1};
					empty_location_en<=1'b1;
					last_state<=BQ1;
					reset_cnt<=1'b1;
					end
			
		    end
			else if(save_en)
			    begin
				occupy_en<=1'b1;
				empty_location_en<=1'b0;
				
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b0;
				if(!rise_fall_end)
					begin
					rise_fall_en_main<=1'b1;
					end
				else
					begin
					rise_fall_en_main<=1'b0;
					end
				if(!rotate_end)
					begin
					rotate_en<=1'b1;
					end
				else
					begin
					rotate_en<=1'b0;
					end
					
				if(S0[6:5]>current_state[6:5])
					begin
					rise_fall_cnt<=(S0[6:5]-current_state[6:5])*RISE_FALL_CNT_A;     //升的高度
					rise_fall_direction<=1'b0;
					end
				else
					begin
					rise_fall_cnt<=(current_state[6:5]-S0[6:5])*RISE_FALL_CNT_A;     //降的高度
					rise_fall_direction<=1'b1;
					end
				if(S0[3:1]>current_state[3:1])
				    begin
				    rotate_cnt<=(S0[3:1]-current_state[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b0;
				    end
				else
				    begin
				    rotate_cnt<=(current_state[3:1]-S0[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b1;
				    end
			    if((!rise_fall_end)|(!rotate_end))
				    begin
					next_state<=BQ1;
					reset_cnt<=1'b0;
				    end
				else
					begin
					next_state<=S0;
					last_state<=BQ1;
					reset_cnt<=1'b1;
					end
			
		        end
			else
				begin
				empty_location_en<=1'b0;
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=BQ1;
				end
		   end
		BQ2:begin
			empty_location_en<=1'b0;
			if(fetch_en)
				begin
				yuyin_end_en<=2'b00;
				accomplish_en<=1'b0;
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=BQ2;
			    	end
			    else
					begin
					last_state<=BQ2;
					next_state<=BQ3;
			    	end
				end
			else if(save_en)
				begin
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b1;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=BQ2;
					occupy_en<=1'b1;
					yuyin_end_en<=2'b00;
					accomplish_en<=1'b0;
			    	end
			    else
					begin
					last_state<=BQ2;
					next_state<=BQ1;
					yuyin_end_en<=2'b01;
					occupy_en<=1'b0;
					accomplish_en<=1'b1;
			    	end
				end
			else
				begin
				yuyin_end_en<=2'b00;
				accomplish_en<=1'b0;
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=BQ2;
				end
		   end
		BQ3:begin
			empty_location_en<=1'b0;
			yuyin_end_en<=2'b00;
			if(fetch_en)
				begin
				occupy_en<=1'b1;
				
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b0;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b1;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=RISE_FALL_CNT_B;     
			    rise_fall_direction<=1'b0;	
				if(!rise_fall_end)
			        begin
					next_state<=BQ3;
			    	end
			    else
					begin
					last_state<=BQ3;
					next_state<=BQ4;
			    	end
				end
			else if(save_en)
				begin
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b0;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b1;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=RISE_FALL_CNT_B;     
			    rise_fall_direction<=1'b1;	
				if(!rise_fall_end)
			        begin
					next_state<=BQ3;
			    	end
			    else
					begin
					last_state<=BQ3;
					next_state<=BQ2;
			    	end
				end
			else
				begin
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=BQ3;
				end
		   end
		BQ4:begin
			empty_location_en<=1'b0;
			yuyin_end_en<=2'b00;
			if(fetch_en)
				begin
				occupy_en<=1'b1;
				
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b1;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=BQ4;
			    	end
			    else
					begin
					last_state<=BQ4;
					next_state<=S3;
			    	end
				end
			else if(save_en)
				begin
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;     //伸缩长度
			    if(!extend_shrink_end)
			        begin
					next_state<=BQ4;
			    	end
			    else
					begin
					last_state<=BQ4;
					next_state<=BQ3;
			    	end
			    end
			else
				begin
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=BQ4;
				end
		   end
		//第二层顺时针第二个房间 
		BW1:begin
		accomplish_en<=1'b0;
		yuyin_end_en<=2'b00;
		    if(fetch_en)
		    begin
				occupy_en<=1'b1;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b0;
				if(!rise_fall_end)
					begin
					rise_fall_en_main<=1'b1;
					end
				else
					begin
					rise_fall_en_main<=1'b0;
					end
				if(!rotate_end)
					begin
					rotate_en<=1'b1;
					end
				else
					begin
					rotate_en<=1'b0;
					end
					
				if(location_coding[6:5]>last_state[6:5])
					begin
					rise_fall_cnt<=(location_coding[6:5]-last_state[6:5])*RISE_FALL_CNT_A;     //升的高度
					rise_fall_direction<=1'b0;
					end
				else
					begin
					rise_fall_cnt<=(last_state[6:5]-location_coding[6:5])*RISE_FALL_CNT_A;     //降的高度
					rise_fall_direction<=1'b1;
					end
				if(location_coding[3:1]>last_state[3:1])
				    begin
				    rotate_cnt<=(location_coding[3:1]-last_state[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b0;
				    end
				else
				    begin
				    rotate_cnt<=(last_state[3:1]-location_coding[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b1;
				    end
			    if((!rise_fall_end)|(!rotate_end))
				    begin
					next_state<=BW1;
					reset_cnt<=1'b0;
				    end
				else
					begin
					next_state<={location_coding[6:1],1'b1};
					empty_location_en<=1'b1;
					last_state<=BW1;
					reset_cnt<=1'b1;
					end
			
		    end
			else if(save_en)
			    begin
				occupy_en<=1'b1;
				empty_location_en<=1'b0;
				
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b0;
				if(!rise_fall_end)
					begin
					rise_fall_en_main<=1'b1;
					end
				else
					begin
					rise_fall_en_main<=1'b0;
					end
				if(!rotate_end)
					begin
					rotate_en<=1'b1;
					end
				else
					begin
					rotate_en<=1'b0;
					end
					
				if(S0[6:5]>current_state[6:5])
					begin
					rise_fall_cnt<=(S0[6:5]-current_state[6:5])*RISE_FALL_CNT_A;     //升的高度
					rise_fall_direction<=1'b0;
					end
				else
					begin
					rise_fall_cnt<=(current_state[6:5]-S0[6:5])*RISE_FALL_CNT_A;     //降的高度
					rise_fall_direction<=1'b1;
					end
				if(S0[3:1]>current_state[3:1])
				    begin
				    rotate_cnt<=(S0[3:1]-current_state[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b0;
				    end
				else
				    begin
				    rotate_cnt<=(current_state[3:1]-S0[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b1;
				    end
			    if((!rise_fall_end)|(!rotate_end))
				    begin
					next_state<=BW1;
					reset_cnt<=1'b0;
				    end
				else
					begin
					next_state<=S0;
					last_state<=BW1;
					reset_cnt<=1'b1;
					end
			
		        end
			else
				begin
				empty_location_en<=1'b0;
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=BW1;
				end
		   end
		BW2:begin
			empty_location_en<=1'b0;
			if(fetch_en)
				begin
				accomplish_en<=1'b0;
				yuyin_end_en<=2'b00;
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=BW2;
			    	end
			    else
					begin
					last_state<=BW2;
					next_state<=BW3;
			    	end
				end
			else if(save_en)
				begin
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b1;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=BW2;
					yuyin_end_en<=2'b00;
					occupy_en<=1'b1;
					accomplish_en<=1'b0;
			    	end
			    else
					begin
					last_state<=BW2;
					next_state<=BW1;
					occupy_en<=1'b0;
					yuyin_end_en<=2'b01;
					accomplish_en<=1'b1;
			    	end
				end
			else
				begin
				accomplish_en<=1'b0;
				occupy_en<=1'b0;
				yuyin_end_en<=2'b00;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=BW2;
				end
		   end
		BW3:begin
			empty_location_en<=1'b0;
			yuyin_end_en<=2'b00;
			if(fetch_en)
				begin
				occupy_en<=1'b1;
				
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b0;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b1;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=RISE_FALL_CNT_B;     
			    rise_fall_direction<=1'b0;	
				if(!rise_fall_end)
			        begin
					next_state<=BW3;
			    	end
			    else
					begin
					last_state<=BW3;
					next_state<=BW4;
			    	end
				end
			else if(save_en)
				begin
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b0;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b1;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=RISE_FALL_CNT_B;     
			    rise_fall_direction<=1'b1;	
				if(!rise_fall_end)
			        begin
					next_state<=BW3;
			    	end
			    else
					begin
					last_state<=BW3;
					next_state<=BW2;
			    	end
				end
			else
				begin
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=BW3;
				end
		   end
		BW4:begin
			empty_location_en<=1'b0;
			yuyin_end_en<=2'b00;
			if(fetch_en)
				begin
				occupy_en<=1'b1;
				
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b1;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=BW4;
			    	end
			    else
					begin
					last_state<=BW4;
					next_state<=S3;
			    	end
				end
			else if(save_en)
				begin
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;     //伸缩长度
			    if(!extend_shrink_end)
			        begin
					next_state<=BW4;
			    	end
			    else
					begin
					last_state<=BW4;
					next_state<=BW3;
			    	end
			    end
			else
				begin
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=BW4;
				end
		   end
		//第二层顺时针第三个房间
		BE1:begin
		accomplish_en<=1'b0;
		yuyin_end_en<=2'b00;
		    if(fetch_en)
		    begin
				occupy_en<=1'b1;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b0;
				if(!rise_fall_end)
					begin
					rise_fall_en_main<=1'b1;
					end
				else
					begin
					rise_fall_en_main<=1'b0;
					end
				if(!rotate_end)
					begin
					rotate_en<=1'b1;
					end
				else
					begin
					rotate_en<=1'b0;
					end
					
				if(location_coding[6:5]>last_state[6:5])
					begin
					rise_fall_cnt<=(location_coding[6:5]-last_state[6:5])*RISE_FALL_CNT_A;     //升的高度
					rise_fall_direction<=1'b0;
					end
				else
					begin
					rise_fall_cnt<=(last_state[6:5]-location_coding[6:5])*RISE_FALL_CNT_A;     //降的高度
					rise_fall_direction<=1'b1;
					end
				if(location_coding[3:1]>last_state[3:1])
				    begin
				    rotate_cnt<=(location_coding[3:1]-last_state[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b0;
				    end
				else
				    begin
				    rotate_cnt<=(last_state[3:1]-location_coding[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b1;
				    end
			    if((!rise_fall_end)|(!rotate_end))
				    begin
					next_state<=BE1;
					reset_cnt<=1'b0;
				    end
				else
					begin
					next_state<={location_coding[6:1],1'b1};
					empty_location_en<=1'b1;
					last_state<=BE1;
					reset_cnt<=1'b1;
					end
			
		    end
			else if(save_en)
			    begin
				occupy_en<=1'b1;
				empty_location_en<=1'b0;
				
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b0;
				if(!rise_fall_end)
					begin
					rise_fall_en_main<=1'b1;
					end
				else
					begin
					rise_fall_en_main<=1'b0;
					end
				if(!rotate_end)
					begin
					rotate_en<=1'b1;
					end
				else
					begin
					rotate_en<=1'b0;
					end
					
				if(S0[6:5]>current_state[6:5])
					begin
					rise_fall_cnt<=(S0[6:5]-current_state[6:5])*RISE_FALL_CNT_A;     //升的高度
					rise_fall_direction<=1'b0;
					end
				else
					begin
					rise_fall_cnt<=(current_state[6:5]-S0[6:5])*RISE_FALL_CNT_A;     //降的高度
					rise_fall_direction<=1'b1;
					end
				if(S0[3:1]>current_state[3:1])
				    begin
				    rotate_cnt<=(S0[3:1]-current_state[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b0;
				    end
				else
				    begin
				    rotate_cnt<=(current_state[3:1]-S0[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b1;
				    end
			    if((!rise_fall_end)|(!rotate_end))
				    begin
					next_state<=BE1;
					reset_cnt<=1'b0;
				    end
				else
					begin
					next_state<=S0;
					last_state<=BE1;
					reset_cnt<=1'b1;
					end
			
		        end
			else
				begin
				empty_location_en<=1'b0;
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=BE1;
				end
		   end
		BE2:begin
			empty_location_en<=1'b0;
			if(fetch_en)
				begin
				accomplish_en<=1'b0;
				yuyin_end_en<=2'b00;
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=BE2;
			    	end
			    else
					begin
					last_state<=BE2;
					next_state<=BE3;
			    	end
				end
			else if(save_en)
				begin
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b1;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=BE2;
					occupy_en<=1'b1;
					accomplish_en<=1'b0;
					yuyin_end_en<=2'b00;
			    	end
			    else
					begin
					yuyin_end_en<=2'b01;
					last_state<=BE2;
					next_state<=BE1;
					occupy_en<=1'b0;
					accomplish_en<=1'b1;
			    	end
				end
			else
				begin
				yuyin_end_en<=2'b00;
				accomplish_en<=1'b0;
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=BE2;
				end
		   end
		BE3:begin
			empty_location_en<=1'b0;
			yuyin_end_en<=2'b00;
			rise_fall_en_main<=1'b0;
			if(fetch_en)
				begin
				occupy_en<=1'b1;
				
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b0;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b1;
				rise_fall_cnt<=RISE_FALL_CNT_B;     
			    rise_fall_direction<=1'b0;	
				if(!rise_fall_end)
			        begin
					next_state<=BE3;
			    	end
			    else
					begin
					last_state<=BE3;
					next_state<=BE4;
			    	end
				end
			else if(save_en)
				begin
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b0;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b1;
				rise_fall_cnt<=RISE_FALL_CNT_B;     
			    rise_fall_direction<=1'b1;	
				if(!rise_fall_end)
			        begin
					next_state<=BE3;
			    	end
			    else
					begin
					last_state<=BE3;
					next_state<=BE2;
			    	end
				end
			else
				begin
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=BE3;
				end
		   end
		BE4:begin
			empty_location_en<=1'b0;
			rise_fall_en_main<=1'b0;
			yuyin_end_en<=2'b00;
			if(fetch_en)
				begin
				occupy_en<=1'b1;
				
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b1;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=BE4;
			    	end
			    else
					begin
					last_state<=BE4;
					next_state<=S3;
			    	end
				end
			else if(save_en)
				begin
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;     //伸缩长度
			    if(!extend_shrink_end)
			        begin
					next_state<=BE4;
			    	end
			    else
					begin
					last_state<=BE4;
					next_state<=BE3;
			    	end
			    end
			else
				begin
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=BE4;
				end
		   end
		//第二层顺时针第四个房间
		BR1:begin
			accomplish_en<=1'b0;
			yuyin_end_en<=2'b00;
		    if(fetch_en)
		    begin
				occupy_en<=1'b1;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b0;
				if(!rise_fall_end)
					begin
					rise_fall_en_main<=1'b1;
					end
				else
					begin
					rise_fall_en_main<=1'b0;
					end
				if(!rotate_end)
					begin
					rotate_en<=1'b1;
					end
				else
					begin
					rotate_en<=1'b0;
					end
					
				if(location_coding[6:5]>last_state[6:5])
					begin
					rise_fall_cnt<=(location_coding[6:5]-last_state[6:5])*RISE_FALL_CNT_A;     //升的高度
					rise_fall_direction<=1'b0;
					end
				else
					begin
					rise_fall_cnt<=(last_state[6:5]-location_coding[6:5])*RISE_FALL_CNT_A;     //降的高度
					rise_fall_direction<=1'b1;
					end
				if(location_coding[3:1]>last_state[3:1])
				    begin
				    rotate_cnt<=(location_coding[3:1]-last_state[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b0;
				    end
				else
				    begin
				    rotate_cnt<=(last_state[3:1]-location_coding[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b1;
				    end
			    if((!rise_fall_end)|(!rotate_end))
				    begin
					next_state<=BR1;
					reset_cnt<=1'b0;
				    end
				else
					begin
					next_state<={location_coding[6:1],1'b1};
					empty_location_en<=1'b1;
					last_state<=BR1;
					reset_cnt<=1'b1;
					end
			
		    end
			else if(save_en)
			    begin
				occupy_en<=1'b1;
				empty_location_en<=1'b0;
				
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b0;
				if(!rise_fall_end)
					begin
					rise_fall_en_main<=1'b1;
					end
				else
					begin
					rise_fall_en_main<=1'b0;
					end
				if(!rotate_end)
					begin
					rotate_en<=1'b1;
					end
				else
					begin
					rotate_en<=1'b0;
					end
					
				if(S0[6:5]>current_state[6:5])
					begin
					rise_fall_cnt<=(S0[6:5]-current_state[6:5])*RISE_FALL_CNT_A;     //升的高度
					rise_fall_direction<=1'b0;
					end
				else
					begin
					rise_fall_cnt<=(current_state[6:5]-S0[6:5])*RISE_FALL_CNT_A;     //降的高度
					rise_fall_direction<=1'b1;
					end
				if(S0[3:1]>current_state[3:1])
				    begin
				    rotate_cnt<=(S0[3:1]-current_state[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b0;
				    end
				else
				    begin
				    rotate_cnt<=(current_state[3:1]-S0[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b1;
				    end
			    if((!rise_fall_end)|(!rotate_end))
				    begin
					next_state<=BR1;
					reset_cnt<=1'b0;
				    end
				else
					begin
					next_state<=S0;
					last_state<=BR1;
					reset_cnt<=1'b1;
					end
			
		        end
			else
				begin
				empty_location_en<=1'b0;
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=BR1;
				end
		   end
		BR2:begin
			rise_fall_en_main<=1'b0;
			empty_location_en<=1'b0;
			if(fetch_en)
				begin
				yuyin_end_en<=2'b00;
				accomplish_en<=1'b0;
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=BR2;
			    	end
			    else
					begin
					last_state<=BR2;
					next_state<=BR3;
			    	end
				end
			else if(save_en)
				begin
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b1;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=BR2;
					occupy_en<=1'b1;
					yuyin_end_en<=2'b00;
					accomplish_en<=1'b0;
			    	end
			    else
					begin
					last_state<=BR2;
					next_state<=BR1;
					yuyin_end_en<=2'b01;
					occupy_en<=1'b0;
					accomplish_en<=1'b1;
			    	end
				end
			else
				begin
				yuyin_end_en<=2'b00;
				accomplish_en<=1'b0;
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=BR2;
				end
		   end
		BR3:begin
			yuyin_end_en<=2'b00;
			empty_location_en<=1'b0;
			rise_fall_en_main<=1'b0;
			if(fetch_en)
				begin
				occupy_en<=1'b1;
				
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b0;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b1;
				rise_fall_cnt<=RISE_FALL_CNT_B;     
			    rise_fall_direction<=1'b0;	
				if(!rise_fall_end)
			        begin
					next_state<=BR3;
			    	end
			    else
					begin
					last_state<=BR3;
					next_state<=BR4;
			    	end
				end
			else if(save_en)
				begin
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b0;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b1;
				rise_fall_cnt<=RISE_FALL_CNT_B;     
			    rise_fall_direction<=1'b1;	
				if(!rise_fall_end)
			        begin
					next_state<=BR3;
			    	end
			    else
					begin
					last_state<=BR3;
					next_state<=BR2;
			    	end
				end
			else
				begin
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=BR3;
				end
		   end
		BR4:begin
			yuyin_end_en<=2'b00;
			empty_location_en<=1'b0;
			rise_fall_en_main<=1'b0;
			if(fetch_en)
				begin
				occupy_en<=1'b1;
				
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b1;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=BR4;
			    	end
			    else
					begin
					last_state<=BR4;
					next_state<=S3;
			    	end
				end
			else if(save_en)
				begin
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;     //伸缩长度
			    if(!extend_shrink_end)
			        begin
					next_state<=BR4;
			    	end
			    else
					begin
					last_state<=BR4;
					next_state<=BR3;
			    	end
			    end
			else
				begin
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=BR4;
				end
		   end
	
//第三层
		//第三层顺时针第一个房间
		CQ1:begin
		accomplish_en<=1'b0;
		yuyin_end_en<=2'b00;
		    if(fetch_en)
		    begin
				occupy_en<=1'b1;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b0;
				if(!rise_fall_end)
					begin
					rise_fall_en_main<=1'b1;
					end
				else
					begin
					rise_fall_en_main<=1'b0;
					end
				if(!rotate_end)
					begin
					rotate_en<=1'b1;
					end
				else
					begin
					rotate_en<=1'b0;
					end
					
				if(location_coding[6:5]>last_state[6:5])
					begin
					rise_fall_cnt<=(location_coding[6:5]-last_state[6:5])*RISE_FALL_CNT_A;     //升的高度
					rise_fall_direction<=1'b0;
					end
				else
					begin
					rise_fall_cnt<=(last_state[6:5]-location_coding[6:5])*RISE_FALL_CNT_A;     //降的高度
					rise_fall_direction<=1'b1;
					end
				if(location_coding[3:1]>last_state[3:1])
				    begin
				    rotate_cnt<=(location_coding[3:1]-last_state[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b0;
				    end
				else
				    begin
				    rotate_cnt<=(last_state[3:1]-location_coding[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b1;
				    end
			    if((!rise_fall_end)|(!rotate_end))
				    begin
					next_state<=CQ1;
					reset_cnt<=1'b0;
				    end
				else
					begin
					next_state<={location_coding[6:1],1'b1};
					empty_location_en<=1'b1;
					last_state<=CQ1;
					reset_cnt<=1'b1;
					end
			
		    end
			else if(save_en)
			    begin
				occupy_en<=1'b1;
				empty_location_en<=1'b0;
				
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b0;
				if(!rise_fall_end)
					begin
					rise_fall_en_main<=1'b1;
					end
				else
					begin
					rise_fall_en_main<=1'b0;
					end
				if(!rotate_end)
					begin
					rotate_en<=1'b1;
					end
				else
					begin
					rotate_en<=1'b0;
					end
					
				if(S0[6:5]>current_state[6:5])
					begin
					rise_fall_cnt<=(S0[6:5]-current_state[6:5])*RISE_FALL_CNT_A;     //升的高度
					rise_fall_direction<=1'b0;
					end
				else
					begin
					rise_fall_cnt<=(current_state[6:5]-S0[6:5])*RISE_FALL_CNT_A;     //降的高度
					rise_fall_direction<=1'b1;
					end
				if(S0[3:1]>current_state[3:1])
				    begin
				    rotate_cnt<=(S0[3:1]-current_state[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b0;
				    end
				else
				    begin
				    rotate_cnt<=(current_state[3:1]-S0[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b1;
				    end
			    if((!rise_fall_end)|(!rotate_end))
				    begin
					next_state<=CQ1;
					reset_cnt<=1'b0;
				    end
				else
					begin
					next_state<=S0;
					last_state<=CQ1;
					reset_cnt<=1'b1;
					end
			
		        end
			else
				begin
				empty_location_en<=1'b0;
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=CQ1;
				end
		   end
		CQ2:begin
			empty_location_en<=1'b0;
			rise_fall_en_main<=1'b0;
			if(fetch_en)
				begin
				yuyin_end_en<=2'b00;
				accomplish_en<=1'b0;
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=CQ2;
			    	end
			    else
					begin
					last_state<=CQ2;
					next_state<=CQ3;
			    	end
				end
			else if(save_en)
				begin
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b1;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=CQ2;
					occupy_en<=1'b1;
					yuyin_end_en<=2'b00;
					accomplish_en<=1'b0;
			    	end
			    else
					begin
					last_state<=CQ2;
					next_state<=CQ1;
					occupy_en<=1'b0;
					yuyin_end_en<=2'b01;
					accomplish_en<=1'b1;
			    	end
				end
			else
				begin
				yuyin_end_en<=2'b00;
				occupy_en<=1'b0;
				accomplish_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=CQ2;
				end
		   end
		CQ3:begin
			yuyin_end_en<=2'b00;
			empty_location_en<=1'b0;
			rise_fall_en_main<=1'b0;
			if(fetch_en)
				begin
				occupy_en<=1'b1;
				
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b0;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b1;
				rise_fall_cnt<=RISE_FALL_CNT_B;     
			    rise_fall_direction<=1'b0;	
				if(!rise_fall_end)
			        begin
					next_state<=CQ3;
			    	end
			    else
					begin
					last_state<=CQ3;
					next_state<=CQ4;
			    	end
				end
			else if(save_en)
				begin
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b0;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b1;
				rise_fall_cnt<=RISE_FALL_CNT_B;     
			    rise_fall_direction<=1'b1;	
				if(!rise_fall_end)
			        begin
					next_state<=CQ3;
			    	end
			    else
					begin
					last_state<=CQ3;
					next_state<=CQ2;
			    	end
				end
			else
				begin
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=CQ3;
				end
		   end
		CQ4:begin
			empty_location_en<=1'b0;
			rise_fall_en_main<=1'b0;
			yuyin_end_en<=2'b00;
			if(fetch_en)
				begin
				occupy_en<=1'b1;
				
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b1;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=CQ4;
			    	end
			    else
					begin
					last_state<=CQ4;
					next_state<=S3;
			    	end
				end
			else if(save_en)
				begin
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;     //伸缩长度
			    if(!extend_shrink_end)
			        begin
					next_state<=CQ4;
			    	end
			    else
					begin
					last_state<=CQ4;
					next_state<=CQ3;
			    	end
			    end
			else
				begin
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=CQ4;
				end
		   end
		//第三层顺时针第二个房间 
		CW1:begin
		accomplish_en<=1'b0;
		yuyin_end_en<=2'b00;
		    if(fetch_en)
		    begin
				occupy_en<=1'b1;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b0;
				if(!rise_fall_end)
					begin
					rise_fall_en_main<=1'b1;
					end
				else
					begin
					rise_fall_en_main<=1'b0;
					end
				if(!rotate_end)
					begin
					rotate_en<=1'b1;
					end
				else
					begin
					rotate_en<=1'b0;
					end
					
				if(location_coding[6:5]>last_state[6:5])
					begin
					rise_fall_cnt<=(location_coding[6:5]-last_state[6:5])*RISE_FALL_CNT_A;     //升的高度
					rise_fall_direction<=1'b0;
					end
				else
					begin
					rise_fall_cnt<=(last_state[6:5]-location_coding[6:5])*RISE_FALL_CNT_A;     //降的高度
					rise_fall_direction<=1'b1;
					end
				if(location_coding[3:1]>last_state[3:1])
				    begin
				    rotate_cnt<=(location_coding[3:1]-last_state[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b0;
				    end
				else
				    begin
				    rotate_cnt<=(last_state[3:1]-location_coding[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b1;
				    end
			    if((!rise_fall_end)|(!rotate_end))
				    begin
					next_state<=CW1;
					reset_cnt<=1'b0;
				    end
				else
					begin
					next_state<={location_coding[6:1],1'b1};
					empty_location_en<=1'b1;
					last_state<=CW1;
					reset_cnt<=1'b1;
					end
			
		    end
			else if(save_en)
			    begin
				occupy_en<=1'b1;
				empty_location_en<=1'b0;
				
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b0;
				if(!rise_fall_end)
					begin
					rise_fall_en_main<=1'b1;
					end
				else
					begin
					rise_fall_en_main<=1'b0;
					end
				if(!rotate_end)
					begin
					rotate_en<=1'b1;
					end
				else
					begin
					rotate_en<=1'b0;
					end
					
				if(S0[6:5]>current_state[6:5])
					begin
					rise_fall_cnt<=(S0[6:5]-current_state[6:5])*RISE_FALL_CNT_A;     //升的高度
					rise_fall_direction<=1'b0;
					end
				else
					begin
					rise_fall_cnt<=(current_state[6:5]-S0[6:5])*RISE_FALL_CNT_A;     //降的高度
					rise_fall_direction<=1'b1;
					end
				if(S0[3:1]>current_state[3:1])
				    begin
				    rotate_cnt<=(S0[3:1]-current_state[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b0;
				    end
				else
				    begin
				    rotate_cnt<=(current_state[3:1]-S0[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b1;
				    end
			    if((!rise_fall_end)|(!rotate_end))
				    begin
					next_state<=CW1;
					reset_cnt<=1'b0;
				    end
				else
					begin
					next_state<=S0;
					last_state<=CW1;
					reset_cnt<=1'b1;
					end
			
		        end
			else
				begin
				empty_location_en<=1'b0;
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=CW1;
				end
		   end
		CW2:begin
			empty_location_en<=1'b0;
			rise_fall_en_main<=1'b0;
			if(fetch_en)
				begin
				yuyin_end_en<=2'b00;
				accomplish_en<=1'b0;
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=CW2;
			    	end
			    else
					begin
					last_state<=CW2;
					next_state<=CW3;
			    	end
				end
			else if(save_en)
				begin
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b1;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=CW2;
					occupy_en<=1'b1;
					yuyin_end_en<=2'b00;
					accomplish_en<=1'b0;
			    	end
			    else
					begin
					last_state<=CW2;
					next_state<=CW1;
					occupy_en<=1'b0;
					yuyin_end_en<=2'b01;
					accomplish_en<=1'b1;
			    	end
				end
			else
				begin
				yuyin_end_en<=2'b00;
				accomplish_en<=1'b0;
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=CW2;
				end
		   end
		CW3:begin
			empty_location_en<=1'b0;
			rise_fall_en_main<=1'b0;
			yuyin_end_en<=2'b00;
			if(fetch_en)
				begin
				occupy_en<=1'b1;
				
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b0;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b1;
				rise_fall_cnt<=RISE_FALL_CNT_B;     
			    rise_fall_direction<=1'b0;	
				if(!rise_fall_end)
			        begin
					next_state<=CW3;
			    	end
			    else
					begin
					last_state<=CW3;
					next_state<=CW4;
			    	end
				end
			else if(save_en)
				begin
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b0;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b1;
				rise_fall_cnt<=RISE_FALL_CNT_B;     
			    rise_fall_direction<=1'b1;	
				if(!rise_fall_end)
			        begin
					next_state<=CW3;
			    	end
			    else
					begin
					last_state<=CW3;
					next_state<=CW2;
			    	end
				end
			else
				begin
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=CW3;
				end
		   end
		CW4:begin
			empty_location_en<=1'b0;
			rise_fall_en_main<=1'b0;
			yuyin_end_en<=2'b00;
			if(fetch_en)
				begin
				occupy_en<=1'b1;
				
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b1;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=CW4;
			    	end
			    else
					begin
					last_state<=CW4;
					next_state<=S3;
			    	end
				end
			else if(save_en)
				begin
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;     //伸缩长度
			    if(!extend_shrink_end)
			        begin
					next_state<=CW4;
			    	end
			    else
					begin
					last_state<=CW4;
					next_state<=CW3;
			    	end
			    end
			else
				begin
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=CW4;
				end
		   end
		//第三层顺时针第三个房间
		CE1:begin
			accomplish_en<=1'b0;
			yuyin_end_en<=2'b00;
		    if(fetch_en)
		    begin
				occupy_en<=1'b1;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b0;
				if(!rise_fall_end)
					begin
					rise_fall_en_main<=1'b1;
					end
				else
					begin
					rise_fall_en_main<=1'b0;
					end
				if(!rotate_end)
					begin
					rotate_en<=1'b1;
					end
				else
					begin
					rotate_en<=1'b0;
					end
					
				if(location_coding[6:5]>last_state[6:5])
					begin
					rise_fall_cnt<=(location_coding[6:5]-last_state[6:5])*RISE_FALL_CNT_A;     //升的高度
					rise_fall_direction<=1'b0;
					end
				else
					begin
					rise_fall_cnt<=(last_state[6:5]-location_coding[6:5])*RISE_FALL_CNT_A;     //降的高度
					rise_fall_direction<=1'b1;
					end
				if(location_coding[3:1]>last_state[3:1])
				    begin
				    rotate_cnt<=(location_coding[3:1]-last_state[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b0;
				    end
				else
				    begin
				    rotate_cnt<=(last_state[3:1]-location_coding[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b1;
				    end
			    if((!rise_fall_end)|(!rotate_end))
				    begin
					next_state<=CE1;
					reset_cnt<=1'b0;
				    end
				else
					begin
					next_state<={location_coding[6:1],1'b1};
					empty_location_en<=1'b1;
					last_state<=CE1;
					reset_cnt<=1'b1;
					end
			
		    end
			else if(save_en)
			    begin
				occupy_en<=1'b1;
				empty_location_en<=1'b0;
				
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b0;
				if(!rise_fall_end)
					begin
					rise_fall_en_main<=1'b1;
					end
				else
					begin
					rise_fall_en_main<=1'b0;
					end
				if(!rotate_end)
					begin
					rotate_en<=1'b1;
					end
				else
					begin
					rotate_en<=1'b0;
					end
					
				if(S0[6:5]>current_state[6:5])
					begin
					rise_fall_cnt<=(S0[6:5]-current_state[6:5])*RISE_FALL_CNT_A;     //升的高度
					rise_fall_direction<=1'b0;
					end
				else
					begin
					rise_fall_cnt<=(current_state[6:5]-S0[6:5])*RISE_FALL_CNT_A;     //降的高度
					rise_fall_direction<=1'b1;
					end
				if(S0[3:1]>current_state[3:1])
				    begin
				    rotate_cnt<=(S0[3:1]-current_state[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b0;
				    end
				else
				    begin
				    rotate_cnt<=(current_state[3:1]-S0[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b1;
				    end
			    if((!rise_fall_end)|(!rotate_end))
				    begin
					next_state<=CE1;
					reset_cnt<=1'b0;
				    end
				else
					begin
					next_state<=S0;
					last_state<=CE1;
					reset_cnt<=1'b1;
					end
			
		        end
			else
				begin
				empty_location_en<=1'b0;
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=CE1;
				end
		   end
		CE2:begin
			empty_location_en<=1'b0;
			rise_fall_en_main<=1'b0;
			if(fetch_en)
				begin
				yuyin_end_en<=2'b00;
				accomplish_en<=1'b0;
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=CE2;
			    	end
			    else
					begin
					last_state<=CE2;
					next_state<=CE3;
			    	end
				end
			else if(save_en)
				begin
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b1;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=CE2;
					occupy_en<=1'b1;
					yuyin_end_en<=2'b00;
					accomplish_en<=1'b0;
			    	end
			    else
					begin
					last_state<=CE2;
					next_state<=CE1;
					occupy_en<=1'b0;
					yuyin_end_en<=2'b01;
					accomplish_en<=1'b1;
			    	end
				end
			else
				begin
				yuyin_end_en<=2'b00;
				accomplish_en<=1'b0;
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=CE2;
				end
		   end
		CE3:begin
			empty_location_en<=1'b0;
			rise_fall_en_main<=1'b0;
			yuyin_end_en<=2'b00;
			if(fetch_en)
				begin
				occupy_en<=1'b1;
				
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b0;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b1;
				rise_fall_cnt<=RISE_FALL_CNT_B;     
			    rise_fall_direction<=1'b0;	
				if(!rise_fall_end)
			        begin
					next_state<=CE3;
			    	end
			    else
					begin
					last_state<=CE3;
					next_state<=CE4;
			    	end
				end
			else if(save_en)
				begin
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b0;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b1;
				rise_fall_cnt<=RISE_FALL_CNT_B;     
			    rise_fall_direction<=1'b1;	
				if(!rise_fall_end)
			        begin
					next_state<=CE3;
			    	end
			    else
					begin
					last_state<=CE3;
					next_state<=CE2;
			    	end
				end
			else
				begin
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=CE3;
				end
		   end
		CE4:begin
			empty_location_en<=1'b0;
			rise_fall_en_main<=1'b0;
			yuyin_end_en<=2'b00;
			if(fetch_en)
				begin
				occupy_en<=1'b1;
				
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b1;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=CE4;
			    	end
			    else
					begin
					last_state<=CE4;
					next_state<=S3;
			    	end
				end
			else if(save_en)
				begin
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;     //伸缩长度
			    if(!extend_shrink_end)
			        begin
					next_state<=CE4;
			    	end
			    else
					begin
					last_state<=CE4;
					next_state<=CE3;
			    	end
			    end
			else
				begin
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=CE4;
				end
		   end
		//第三层顺时针第四个房间
		CR1:begin
		accomplish_en<=1'b0;
		yuyin_end_en<=2'b00;
		    if(fetch_en)
		    begin
				occupy_en<=1'b1;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b0;
				if(!rise_fall_end)
					begin
					rise_fall_en_main<=1'b1;
					end
				else
					begin
					rise_fall_en_main<=1'b0;
					end
				if(!rotate_end)
					begin
					rotate_en<=1'b1;
					end
				else
					begin
					rotate_en<=1'b0;
					end
					
				if(location_coding[6:5]>last_state[6:5])
					begin
					rise_fall_cnt<=(location_coding[6:5]-last_state[6:5])*RISE_FALL_CNT_A;     //升的高度
					rise_fall_direction<=1'b0;
					end
				else
					begin
					rise_fall_cnt<=(last_state[6:5]-location_coding[6:5])*RISE_FALL_CNT_A;     //降的高度
					rise_fall_direction<=1'b1;
					end
				if(location_coding[3:1]>last_state[3:1])
				    begin
				    rotate_cnt<=(location_coding[3:1]-last_state[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b0;
				    end
				else
				    begin
				    rotate_cnt<=(last_state[3:1]-location_coding[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b1;
				    end
			    if((!rise_fall_end)|(!rotate_end))
				    begin
					next_state<=CR1;
					reset_cnt<=1'b0;
				    end
				else
					begin
					next_state<={location_coding[6:1],1'b1};
					empty_location_en<=1'b1;
					last_state<=CR1;
					reset_cnt<=1'b1;
					end
			
		    end
			else if(save_en)
			    begin
				occupy_en<=1'b1;
				empty_location_en<=1'b0;
				
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b0;
				if(!rise_fall_end)
					begin
					rise_fall_en_main<=1'b1;
					end
				else
					begin
					rise_fall_en_main<=1'b0;
					end
				if(!rotate_end)
					begin
					rotate_en<=1'b1;
					end
				else
					begin
					rotate_en<=1'b0;
					end
					
				if(S0[6:5]>current_state[6:5])
					begin
					rise_fall_cnt<=(S0[6:5]-current_state[6:5])*RISE_FALL_CNT_A;     //升的高度
					rise_fall_direction<=1'b0;
					end
				else
					begin
					rise_fall_cnt<=(current_state[6:5]-S0[6:5])*RISE_FALL_CNT_A;     //降的高度
					rise_fall_direction<=1'b1;
					end
				if(S0[3:1]>current_state[3:1])
				    begin
				    rotate_cnt<=(S0[3:1]-current_state[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b0;
				    end
				else
				    begin
				    rotate_cnt<=(current_state[3:1]-S0[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b1;
				    end
			    if((!rise_fall_end)|(!rotate_end))
				    begin
					next_state<=CR1;
					reset_cnt<=1'b0;
				    end
				else
					begin
					next_state<=S0;
					last_state<=CR1;
					reset_cnt<=1'b1;
					end
			
		        end
			else
				begin
				empty_location_en<=1'b0;
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=CR1;
				end
		   end
		CR2:begin
			empty_location_en<=1'b0;
			rise_fall_en_main<=1'b0;
			if(fetch_en)
				begin
				yuyin_end_en<=2'b00;
				accomplish_en<=1'b0;
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=CR2;
			    	end
			    else
					begin
					last_state<=CR2;
					next_state<=CR3;
			    	end
				end
			else if(save_en)
				begin
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b1;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=CR2;
					occupy_en<=1'b1;
					yuyin_end_en<=2'b00;
					accomplish_en<=1'b0;
			    	end
			    else
					begin
					last_state<=CR2;
					next_state<=CR1;
					occupy_en<=1'b0;
					yuyin_end_en<=2'b01;
					accomplish_en<=1'b1;
			    	end
				end
			else
				begin
				yuyin_end_en<=2'b00;
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				accomplish_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=CR2;
				end
		   end
		CR3:begin
			empty_location_en<=1'b0;
			rise_fall_en_main<=1'b0;
			yuyin_end_en<=2'b00;
			if(fetch_en)
				begin
				occupy_en<=1'b1;
				
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b0;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b1;
				rise_fall_cnt<=RISE_FALL_CNT_B;     
			    rise_fall_direction<=1'b0;	
				if(!rise_fall_end)
			        begin
					next_state<=CR3;
			    	end
			    else
					begin
					last_state<=CR3;
					next_state<=CR4;
			    	end
				end
			else if(save_en)
				begin
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b0;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b1;
				rise_fall_cnt<=RISE_FALL_CNT_B;     
			    rise_fall_direction<=1'b1;	
				if(!rise_fall_end)
			        begin
					next_state<=CR3;
			    	end
			    else
					begin
					last_state<=CR3;
					next_state<=CR2;
			    	end
				end
			else
				begin
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=CR3;
				end
		   end
		CR4:begin
			empty_location_en<=1'b0;
			rise_fall_en_main<=1'b0;
			yuyin_end_en<=2'b00;
			if(fetch_en)
				begin
				occupy_en<=1'b1;
				
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b1;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=CR4;
			    	end
			    else
					begin
					last_state<=CR4;
					next_state<=S3;
			    	end
				end
			else if(save_en)
				begin
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;     //伸缩长度
			    if(!extend_shrink_end)
			        begin
					next_state<=CR4;
			    	end
			    else
					begin
					last_state<=CR4;
					next_state<=CR3;
			    	end
			    end
			else
				begin
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=CR4;
				end
		   end
		
//第四层
		//第四层顺时针第一个房间
		DQ1:begin
		yuyin_end_en<=2'b00;
		accomplish_en<=1'b0;
		    if(fetch_en)
		    begin
				occupy_en<=1'b1;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b0;
				if(!rise_fall_end)
					begin
					rise_fall_en_main<=1'b1;
					end
				else
					begin
					rise_fall_en_main<=1'b0;
					end
				if(!rotate_end)
					begin
					rotate_en<=1'b1;
					end
				else
					begin
					rotate_en<=1'b0;
					end
					
				if(location_coding[6:5]>last_state[6:5])
					begin
					rise_fall_cnt<=(location_coding[6:5]-last_state[6:5])*RISE_FALL_CNT_A;     //升的高度
					rise_fall_direction<=1'b0;
					end
				else
					begin
					rise_fall_cnt<=(last_state[6:5]-location_coding[6:5])*RISE_FALL_CNT_A;     //降的高度
					rise_fall_direction<=1'b1;
					end
				if(location_coding[3:1]>last_state[3:1])
				    begin
				    rotate_cnt<=(location_coding[3:1]-last_state[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b0;
				    end
				else
				    begin
				    rotate_cnt<=(last_state[3:1]-location_coding[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b1;
				    end
			    if((!rise_fall_end)|(!rotate_end))
				    begin
					next_state<=DQ1;
					reset_cnt<=1'b0;
				    end
				else
					begin
					next_state<={location_coding[6:1],1'b1};
					empty_location_en<=1'b1;
					last_state<=DQ1;
					reset_cnt<=1'b1;
					end
			
		    end
			else if(save_en)
			    begin
				occupy_en<=1'b1;
				empty_location_en<=1'b0;
				
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b0;
				if(!rise_fall_end)
					begin
					rise_fall_en_main<=1'b1;
					end
				else
					begin
					rise_fall_en_main<=1'b0;
					end
				if(!rotate_end)
					begin
					rotate_en<=1'b1;
					end
				else
					begin
					rotate_en<=1'b0;
					end
					
				if(S0[6:5]>current_state[6:5])
					begin
					rise_fall_cnt<=(S0[6:5]-current_state[6:5])*RISE_FALL_CNT_A;     //升的高度
					rise_fall_direction<=1'b0;
					end
				else
					begin
					rise_fall_cnt<=(current_state[6:5]-S0[6:5])*RISE_FALL_CNT_A;     //降的高度
					rise_fall_direction<=1'b1;
					end
				if(S0[3:1]>current_state[3:1])
				    begin
				    rotate_cnt<=(S0[3:1]-current_state[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b0;
				    end
				else
				    begin
				    rotate_cnt<=(current_state[3:1]-S0[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b1;
				    end
			    if((!rise_fall_end)|(!rotate_end))
				    begin
					next_state<=DQ1;
					reset_cnt<=1'b0;
				    end
				else
					begin
					next_state<=S0;
					last_state<=DQ1;
					reset_cnt<=1'b1;
					end
			
		        end
			else
				begin
				empty_location_en<=1'b0;
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=DQ1;
				end
		   end
		DQ2:begin
			empty_location_en<=1'b0;
			rise_fall_en_main<=1'b0;
			if(fetch_en)
				begin
				yuyin_end_en<=2'b00;
				accomplish_en<=1'b0;
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=DQ2;
			    	end
			    else
					begin
					last_state<=DQ2;
					next_state<=DQ3;
			    	end
				end
			else if(save_en)
				begin
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b1;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=DQ2;
					occupy_en<=1'b1;
					yuyin_end_en<=2'b00;
					accomplish_en<=1'b0;
			    	end
			    else
					begin
					last_state<=DQ2;
					next_state<=DQ1;
					occupy_en<=1'b0;
					yuyin_end_en<=2'b01;
					accomplish_en<=1'b1;
			    	end
				end
			else
				begin
				yuyin_end_en<=2'b00;
				accomplish_en<=1'b0;
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=DQ2;
				end
		   end
		DQ3:begin
			yuyin_end_en<=2'b00;
			empty_location_en<=1'b0;
			rise_fall_en_main<=1'b0;
			if(fetch_en)
				begin
				occupy_en<=1'b1;
				
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b0;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b1;
				rise_fall_cnt<=RISE_FALL_CNT_B;     
			    rise_fall_direction<=1'b0;	
				if(!rise_fall_end)
			        begin
					next_state<=DQ3;
			    	end
			    else
					begin
					last_state<=DQ3;
					next_state<=DQ4;
			    	end
				end
			else if(save_en)
				begin
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b0;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b1;
				rise_fall_cnt<=RISE_FALL_CNT_B;     
			    rise_fall_direction<=1'b1;	
				if(!rise_fall_end)
			        begin
					next_state<=DQ3;
			    	end
			    else
					begin
					last_state<=DQ3;
					next_state<=DQ2;
			    	end
				end
			else
				begin
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=DQ3;
				end
		   end
		DQ4:begin
			yuyin_end_en<=2'b00;
			empty_location_en<=1'b0;
			rise_fall_en_main<=1'b0;
			if(fetch_en)
				begin
				occupy_en<=1'b1;
				
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b1;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=DQ4;
			    	end
			    else
					begin
					last_state<=DQ4;
					next_state<=S3;
			    	end
				end
			else if(save_en)
				begin
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;     //伸缩长度
			    if(!extend_shrink_end)
			        begin
					next_state<=DQ4;
			    	end
			    else
					begin
					last_state<=DQ4;
					next_state<=DQ3;
			    	end
			    end
			else
				begin
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=DQ4;
				end
		   end
		//第四层顺时针第二个房间
		DW1:begin
		accomplish_en<=1'b0;
		yuyin_end_en<=2'b00;
		    if(fetch_en)
		    begin
				occupy_en<=1'b1;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b0;
				if(!rise_fall_end)
					begin
					rise_fall_en_main<=1'b1;
					end
				else
					begin
					rise_fall_en_main<=1'b0;
					end
				if(!rotate_end)
					begin
					rotate_en<=1'b1;
					end
				else
					begin
					rotate_en<=1'b0;
					end
					
				if(location_coding[6:5]>last_state[6:5])
					begin
					rise_fall_cnt<=(location_coding[6:5]-last_state[6:5])*RISE_FALL_CNT_A;     //升的高度
					rise_fall_direction<=1'b0;
					end
				else
					begin
					rise_fall_cnt<=(last_state[6:5]-location_coding[6:5])*RISE_FALL_CNT_A;     //降的高度
					rise_fall_direction<=1'b1;
					end
				if(location_coding[3:1]>last_state[3:1])
				    begin
				    rotate_cnt<=(location_coding[3:1]-last_state[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b0;
				    end
				else
				    begin
				    rotate_cnt<=(last_state[3:1]-location_coding[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b1;
				    end
			    if((!rise_fall_end)|(!rotate_end))
				    begin
					next_state<=DW1;
					reset_cnt<=1'b0;
				    end
				else
					begin
					next_state<={location_coding[6:1],1'b1};
					empty_location_en<=1'b1;
					last_state<=DW1;
					reset_cnt<=1'b1;
					end
			
		    end
			else if(save_en)
			    begin
				occupy_en<=1'b1;
				empty_location_en<=1'b0;
				
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b0;
				if(!rise_fall_end)
					begin
					rise_fall_en_main<=1'b1;
					end
				else
					begin
					rise_fall_en_main<=1'b0;
					end
				if(!rotate_end)
					begin
					rotate_en<=1'b1;
					end
				else
					begin
					rotate_en<=1'b0;
					end
					
				if(S0[6:5]>current_state[6:5])
					begin
					rise_fall_cnt<=(S0[6:5]-current_state[6:5])*RISE_FALL_CNT_A;     //升的高度
					rise_fall_direction<=1'b0;
					end
				else
					begin
					rise_fall_cnt<=(current_state[6:5]-S0[6:5])*RISE_FALL_CNT_A;     //降的高度
					rise_fall_direction<=1'b1;
					end
				if(S0[3:1]>current_state[3:1])
				    begin
				    rotate_cnt<=(S0[3:1]-current_state[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b0;
				    end
				else
				    begin
				    rotate_cnt<=(current_state[3:1]-S0[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b1;
				    end
			    if((!rise_fall_end)|(!rotate_end))
				    begin
					next_state<=DW1;
					reset_cnt<=1'b0;
				    end
				else
					begin
					next_state<=S0;
					last_state<=DW1;
					reset_cnt<=1'b1;
					end
			
		        end
			else
				begin
				empty_location_en<=1'b0;
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=DW1;
				end
		   end
		DW2:begin
			empty_location_en<=1'b0;
			rise_fall_en_main<=1'b0;
			if(fetch_en)
				begin
				yuyin_end_en<=2'b00;
				accomplish_en<=1'b0;
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=DW2;
			    	end
			    else
					begin
					last_state<=DW2;
					next_state<=DW3;
			    	end
				end
			else if(save_en)
				begin
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b1;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=DW2;
					occupy_en<=1'b1;
					yuyin_end_en<=2'b00;
					accomplish_en<=1'b0;
			    	end
			    else
					begin
					last_state<=DW2;
					next_state<=DW1;
					yuyin_end_en<=2'b01;
					occupy_en<=1'b0;
					accomplish_en<=1'b1;
			    	end
				end
			else
				begin
				accomplish_en<=1'b0;
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				yuyin_end_en<=2'b00;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=DW2;
				end
		   end
		DW3:begin
			empty_location_en<=1'b0;
			rise_fall_en_main<=1'b0;
			yuyin_end_en<=2'b00;
			if(fetch_en)
				begin
				occupy_en<=1'b1;
				
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b0;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b1;
				rise_fall_cnt<=RISE_FALL_CNT_B;     
			    rise_fall_direction<=1'b0;	
				if(!rise_fall_end)
			        begin
					next_state<=DW3;
			    	end
			    else
					begin
					last_state<=DW3;
					next_state<=DW4;
			    	end
				end
			else if(save_en)
				begin
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b0;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b1;
				rise_fall_cnt<=RISE_FALL_CNT_B;     
			    rise_fall_direction<=1'b1;	
				if(!rise_fall_end)
			        begin
					next_state<=DW3;
			    	end
			    else
					begin
					last_state<=DW3;
					next_state<=DW2;
			    	end
				end
			else
				begin
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=DW3;
				end
		   end
		DW4:begin
			empty_location_en<=1'b0;
			rise_fall_en_main<=1'b0;
			yuyin_end_en<=2'b00;
			if(fetch_en)
				begin
				occupy_en<=1'b1;
				
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b1;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=DW4;
			    	end
			    else
					begin
					last_state<=DW4;
					next_state<=S3;
			    	end
				end
			else if(save_en)
				begin
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;     //伸缩长度
			    if(!extend_shrink_end)
			        begin
					next_state<=DW4;
			    	end
			    else
					begin
					last_state<=DW4;
					next_state<=DW3;
			    	end
			    end
			else
				begin
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=DW4;
				end
		   end
		//第四层顺时针第三个房间
		DE1:begin
		accomplish_en<=1'b0;
		yuyin_end_en<=2'b00;
		    if(fetch_en)
		    begin
				occupy_en<=1'b1;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b0;
				if(!rise_fall_end)
					begin
					rise_fall_en_main<=1'b1;
					end
				else
					begin
					rise_fall_en_main<=1'b0;
					end
				if(!rotate_end)
					begin
					rotate_en<=1'b1;
					end
				else
					begin
					rotate_en<=1'b0;
					end
					
				if(location_coding[6:5]>last_state[6:5])
					begin
					rise_fall_cnt<=(location_coding[6:5]-last_state[6:5])*RISE_FALL_CNT_A;     //升的高度
					rise_fall_direction<=1'b0;
					end
				else
					begin
					rise_fall_cnt<=(last_state[6:5]-location_coding[6:5])*RISE_FALL_CNT_A;     //降的高度
					rise_fall_direction<=1'b1;
					end
				if(location_coding[3:1]>last_state[3:1])
				    begin
				    rotate_cnt<=(location_coding[3:1]-last_state[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b0;
				    end
				else
				    begin
				    rotate_cnt<=(last_state[3:1]-location_coding[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b1;
				    end
			    if((!rise_fall_end)|(!rotate_end))
				    begin
					next_state<=DE1;
					reset_cnt<=1'b0;
				    end
				else
					begin
					next_state<={location_coding[6:1],1'b1};
					empty_location_en<=1'b1;
					last_state<=DE1;
					reset_cnt<=1'b1;
					end
			
		    end
			else if(save_en)
			    begin
				occupy_en<=1'b1;
				empty_location_en<=1'b0;
				
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b0;
				if(!rise_fall_end)
					begin
					rise_fall_en_main<=1'b1;
					end
				else
					begin
					rise_fall_en_main<=1'b0;
					end
				if(!rotate_end)
					begin
					rotate_en<=1'b1;
					end
				else
					begin
					rotate_en<=1'b0;
					end
					
				if(S0[6:5]>current_state[6:5])
					begin
					rise_fall_cnt<=(S0[6:5]-current_state[6:5])*RISE_FALL_CNT_A;     //升的高度
					rise_fall_direction<=1'b0;
					end
				else
					begin
					rise_fall_cnt<=(current_state[6:5]-S0[6:5])*RISE_FALL_CNT_A;     //降的高度
					rise_fall_direction<=1'b1;
					end
				if(S0[3:1]>current_state[3:1])
				    begin
				    rotate_cnt<=(S0[3:1]-current_state[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b0;
				    end
				else
				    begin
				    rotate_cnt<=(current_state[3:1]-S0[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b1;
				    end
			    if((!rise_fall_end)|(!rotate_end))
				    begin
					next_state<=DE1;
					reset_cnt<=1'b0;
				    end
				else
					begin
					next_state<=S0;
					last_state<=DE1;
					reset_cnt<=1'b1;
					end
			
		        end
			else
				begin
				empty_location_en<=1'b0;
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=DE1;
				end
		   end
		DE2:begin
			empty_location_en<=1'b0;
			rise_fall_en_main<=1'b0;
			if(fetch_en)
				begin
				yuyin_end_en<=2'b00;
				accomplish_en<=1'b0;
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=DE2;
			    	end
			    else
					begin
					last_state<=DE2;
					next_state<=DE3;
			    	end
				end
			else if(save_en)
				begin
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b1;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=DE2;
					accomplish_en<=1'b0;
					yuyin_end_en<=2'b00;
					occupy_en<=1'b1;
			    	end
			    else
					begin
					last_state<=DE2;
					next_state<=DE1;
					occupy_en<=1'b0;
					yuyin_end_en<=2'b01;
					accomplish_en<=1'b1;
			    	end
				end
			else
				begin
				yuyin_end_en<=2'b00;
				accomplish_en<=1'b0;
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=DE2;
				end
		   end
		DE3:begin
			yuyin_end_en<=2'b00;
			empty_location_en<=1'b0;
			rise_fall_en_main<=1'b0;
			if(fetch_en)
				begin
				occupy_en<=1'b1;
				
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b0;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b1;
				rise_fall_cnt<=RISE_FALL_CNT_B;     
			    rise_fall_direction<=1'b0;	
				if(!rise_fall_end)
			        begin
					next_state<=DE3;
			    	end
			    else
					begin
					last_state<=DE3;
					next_state<=DE4;
			    	end
				end
			else if(save_en)
				begin
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b0;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b1;
				rise_fall_cnt<=RISE_FALL_CNT_B;     
			    rise_fall_direction<=1'b1;	
				if(!rise_fall_end)
			        begin
					next_state<=DE3;
			    	end
			    else
					begin
					last_state<=DE3;
					next_state<=DE2;
			    	end
				end
			else
				begin
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=DE3;
				end
		   end
		DE4:begin
			yuyin_end_en<=2'b00;
			empty_location_en<=1'b0;
			rise_fall_en_main<=1'b0;
			if(fetch_en)
				begin
				occupy_en<=1'b1;
				
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b1;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=DE4;
			    	end
			    else
					begin
					last_state<=DE4;
					next_state<=S3;
			    	end
				end
			else if(save_en)
				begin
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;     //伸缩长度
			    if(!extend_shrink_end)
			        begin
					next_state<=DE4;
			    	end
			    else
					begin
					last_state<=DE4;
					next_state<=DE3;
			    	end
			    end
			else
				begin
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=DE4;
				end
		   end
		//第四层顺时针第四个房间
		DR1:begin
			yuyin_end_en<=2'b00;
			accomplish_en<=1'b0;
		    if(fetch_en)
		    begin
				occupy_en<=1'b1;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b0;
				if(!rise_fall_end)
					begin
					rise_fall_en_main<=1'b1;
					end
				else
					begin
					rise_fall_en_main<=1'b0;
					end
				if(!rotate_end)
					begin
					rotate_en<=1'b1;
					end
				else
					begin
					rotate_en<=1'b0;
					end
					
				if(location_coding[6:5]>last_state[6:5])
					begin
					rise_fall_cnt<=(location_coding[6:5]-last_state[6:5])*RISE_FALL_CNT_A;     //升的高度
					rise_fall_direction<=1'b0;
					end
				else
					begin
					rise_fall_cnt<=(last_state[6:5]-location_coding[6:5])*RISE_FALL_CNT_A;     //降的高度
					rise_fall_direction<=1'b1;
					end
				if(location_coding[3:1]>last_state[3:1])
				    begin
				    rotate_cnt<=(location_coding[3:1]-last_state[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b0;
				    end
				else
				    begin
				    rotate_cnt<=(last_state[3:1]-location_coding[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b1;
				    end
			    if((!rise_fall_end)|(!rotate_end))
				    begin
					next_state<=DR1;
					reset_cnt<=1'b0;
				    end
				else
					begin
					next_state<={location_coding[6:1],1'b1};
					empty_location_en<=1'b1;
					last_state<=DR1;
					reset_cnt<=1'b1;
					end
			
		    end
			else if(save_en)
			    begin
				occupy_en<=1'b1;
				empty_location_en<=1'b0;
				
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b0;
				if(!rise_fall_end)
					begin
					rise_fall_en_main<=1'b1;
					end
				else
					begin
					rise_fall_en_main<=1'b0;
					end
				if(!rotate_end)
					begin
					rotate_en<=1'b1;
					end
				else
					begin
					rotate_en<=1'b0;
					end
					
				if(S0[6:5]>current_state[6:5])
					begin
					rise_fall_cnt<=(S0[6:5]-current_state[6:5])*RISE_FALL_CNT_A;     //升的高度
					rise_fall_direction<=1'b0;
					end
				else
					begin
					rise_fall_cnt<=(current_state[6:5]-S0[6:5])*RISE_FALL_CNT_A;     //降的高度
					rise_fall_direction<=1'b1;
					end
				if(S0[3:1]>current_state[3:1])
				    begin
				    rotate_cnt<=(S0[3:1]-current_state[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b0;
				    end
				else
				    begin
				    rotate_cnt<=(current_state[3:1]-S0[3:1])*ROTATE_CNT_A;
					rotate_direction<=1'b1;
				    end
			    if((!rise_fall_end)|(!rotate_end))
				    begin
					next_state<=DR1;
					reset_cnt<=1'b0;
				    end
				else
					begin
					next_state<=S0;
					last_state<=DR1;
					reset_cnt<=1'b1;
					end
			
		        end
			else
				begin
				empty_location_en<=1'b0;
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_en_main<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=DR1;
				end
		   end
		DR2:begin
			empty_location_en<=1'b0;
			rise_fall_en_main<=1'b0;
			if(fetch_en)
				begin
				yuyin_end_en<=2'b00;
				accomplish_en<=1'b0;
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=DR2;
			    	end
			    else
					begin
					last_state<=DR2;
					next_state<=DR3;
			    	end
				end
			else if(save_en)
				begin
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b1;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=DR2;
					occupy_en<=1'b1;
					yuyin_end_en<=2'b00;
					accomplish_en<=1'b0;
			    	end
			    else
					begin
					last_state<=DR2;
					next_state<=DR1;
					yuyin_end_en<=2'b01;
					occupy_en<=1'b0;
					accomplish_en<=1'b1;
			    	end
				end
			else
				begin
				yuyin_end_en<=2'b00;
				accomplish_en<=1'b0;
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=DR2;
				end
		   end
		DR3:begin
			empty_location_en<=1'b0;
			rise_fall_en_main<=1'b0;
			yuyin_end_en<=2'b00;
			if(fetch_en)
				begin
				occupy_en<=1'b1;
				
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b0;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b1;
				rise_fall_cnt<=RISE_FALL_CNT_B;     
			    rise_fall_direction<=1'b0;	
				if(!rise_fall_end)
			        begin
					next_state<=DR3;
			    	end
			    else
					begin
					last_state<=DR3;
					next_state<=DR4;
			    	end
				end
			else if(save_en)
				begin
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b0;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=32'd0;
				rise_fall_en<=1'b1;
				rise_fall_cnt<=RISE_FALL_CNT_B;     
			    rise_fall_direction<=1'b1;	
				if(!rise_fall_end)
			        begin
					next_state<=DR3;
			    	end
			    else
					begin
					last_state<=DR3;
					next_state<=DR2;
			    	end
				end
			else
				begin
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=DR3;
				end
		   end
		DR4:begin
			empty_location_en<=1'b0;
			rise_fall_en_main<=1'b0;
			yuyin_end_en<=2'b00;
			if(fetch_en)
				begin
				occupy_en<=1'b1;
				
				rotate_en<=1'b0;
				rotate_cnt<=32'd0;
				rotate_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b1;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;	
				if(!extend_shrink_end)
			        begin
					next_state<=DR4;
			    	end
			    else
					begin
					last_state<=DR4;
					next_state<=S3;
			    	end
				end
			else if(save_en)
				begin
				occupy_en<=1'b1;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				extend_shrink_en<=1'b1;
				extend_shrink_direction<=1'b0;
				extend_shrink_cnt<=EXTEND_SHRINK_CNT_A;     //伸缩长度
			    if(!extend_shrink_end)
			        begin
					next_state<=DR4;
			    	end
			    else
					begin
					last_state<=DR4;
					next_state<=DR3;
			    	end
			    end
			else
				begin
				occupy_en<=1'b0;
				rotate_en<=1'b0;
				rotate_direction<=1'b0;
				rotate_cnt<=32'd0;
				extend_shrink_en<=1'b0;
				extend_shrink_cnt<=32'd0;
				extend_shrink_direction<=1'b0;
				rise_fall_en<=1'b0;
				rise_fall_cnt<=32'd0;     
			    rise_fall_direction<=1'b0;
				next_state<=DR4;
				end
		   end
		
		
		   endcase
		end
	end
	
	
////////////////////////////////////////////////////////////计数器模块//////////////////////////	
	always@(posedge clk or negedge rst_n)
	begin
	if(!rst_n)
		begin
		extend_shrink_end<=1'b0;
		cnt_a<=32'd0;
		end
	else if(extend_shrink_en)
		begin
		if(cnt_a==extend_shrink_cnt)
			begin
			extend_shrink_end<=1'b1;
			cnt_a<=cnt_a;
			end
		else
		    begin
			cnt_a<=cnt_a+1'b1;
			extend_shrink_end<=1'b0;
			end
		end
	else
		begin
		extend_shrink_end<=2'b0;
		cnt_a<=32'd0;
		end
	end
	
	always@(posedge clk or negedge rst_n)
	begin
	if(!rst_n)
		begin
		rise_fall_end<=1'b0;
		cnt_b<=32'd0;
		end
	else if(rise_fall_en|rise_fall_en_main)
		begin
		if(cnt_b==rise_fall_cnt)
			begin
			rise_fall_end<=1'b1;
			cnt_b<=cnt_b;
			end
		else
		    begin
			cnt_b<=cnt_b+1'b1;
			rise_fall_end<=1'b0;
			end
		end
	else if(!reset_cnt)
		begin
		rise_fall_end<=rise_fall_end;
		cnt_b<=cnt_b;
		end
	else 
		begin
		rise_fall_end<=1'b0;
		cnt_b<=32'd0;
		end
	end
	
	always@(posedge clk or negedge rst_n)
	begin
	if(!rst_n)
		begin
		rotate_end<=1'b0;
		cnt_c<=32'd0;
		end
	else if(rotate_en)
		begin
		if(cnt_c==rotate_cnt)
			begin
			rotate_end<=1'b1;
			cnt_c<=cnt_c;
			end
		else
		    begin
			cnt_c<=cnt_c+1'b1;
			rotate_end<=1'b0;
			end
		end
	else if(!reset_cnt)
		begin
		rotate_end<=rotate_end;
		cnt_c<=cnt_c;
		end
	else
		begin
		rotate_end<=1'b0;
		cnt_c<=32'd0;
		end
	end
	
endmodule
